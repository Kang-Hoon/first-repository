module f_not (A,Q);
    input A;
    output Q;
    assign Q    = !A ; 
endmodule